////////////////////////////////////////////////////////////////////////////////
// SubModule 10M08SAE144
// Created   01/02/2015 23:25:02
////////////////////////////////////////////////////////////////////////////////

module 10M08SAE144 (Thermal, GND__142, GND__137, GND__133, GND__125, GND__116, GND__104, GND__95, GND__83, GND__68, GND__63, GND__53, GND__42, REFGND__4, ANAIN1__3, ADC_VREF__5, INPUT_ONLY_8_129/NCONFIG, IO_8_138/CONF_DONE/DIFFIO_RX_T24N, IO_8_136/NSTATUS/DIFFIO_RX_T24P, IO_8_134/CRC_ERROR/DIFFIO_RX_T22N, IO_8_126/BOOT_SEL, IO_8_122/DEV_OE/DIFFIO_RX_T18P, IO_8_121/DEV_CLRN/DIFFIO_RX_T16N, IO_1B_20/TDO/DIFFIO_RX_L12P, IO_1B_19/TDI/DIFFIO_RX_L12N, IO_1B_18/TCK/DIFFIO_RX_L11P, IO_1B_16/TMS/DIFFIO_RX_L11N, IO_1B_15/JTAGEN/DIFFIO_RX_L9P, IO_8_123/VREFB8N0, IO_7_112/VREFB7N0, IO_6_97/VREFB6N0, IO_5_80/VREFB5N0, IO_4_61/VREFB4N0, IO_3_48/VREFB3N0, IO_2_30/VREFB2N0, IO_1B_17/VREFB1N0, IO_6_98/DPCLK2/DIFFIO_RX_R26N, IO_6_96/DPCLK3/DIFFIO_RX_R26P, IO_6_91/CLK3N/DIFFIO_RX_R16N, IO_6_90/CLK3P/DIFFIO_RX_R16P, IO_6_89/CLK2N/DIFFIO_RX_R14N, IO_6_88/CLK2P/DIFFIO_RX_R14P, IO_2_29/CLK1P/DIFFIO_RX_L20P, IO_2_28/CLK1N/DIFFIO_RX_L20N, IO_2_27/CLK0P/DIFFIO_RX_L18P, IO_2_26/CLK0N/DIFFIO_RX_L18N, IO_8_120/DIFFIO_RX_T16P, IO_8_141/DIFFIO_RX_T26N, IO_8_140/DIFFIO_RX_T26P, IO_8_135/DIFFIO_RX_T23N, IO_8_132/DIFFIO_RX_T22P, IO_8_131/DIFFIO_RX_T20N, IO_8_130/DIFFIO_RX_T20P, IO_8_127/DIFFIO_RX_T19N, IO_8_124/DIFFIO_RX_T19P, IO_7_119/DIFFIO_RX_T10N, IO_7_118/DIFFIO_RX_T10P, IO_7_114/DIFFIO_RX_T6P, IO_7_113/DIFFIO_RX_T4N, IO_7_111/DIFFIO_RX_T1N, IO_7_110/DIFFIO_RX_T1P, IO_6_106/DIFFIO_RX_R33N, IO_6_105/DIFFIO_RX_R33P, IO_6_102/DIFFIO_RX_R28N, IO_6_101/DIFFIO_RX_R27N, IO_6_100/DIFFIO_RX_R28P, IO_6_99/DIFFIO_RX_R27P, IO_6_93/DIFFIO_RX_R18N, IO_6_92/DIFFIO_RX_R18P, IO_5_86/DIFFIO_RX_R11N, IO_5_87/DIFFIO_RX_R10N, IO_5_84/DIFFIO_RX_R11P, IO_5_85/DIFFIO_RX_R10P, IO_5_81/DIFFIO_RX_R7N, IO_5_78, IO_5_79/DIFFIO_RX_R7P, IO_5_76/DIFFIO_RX_R2N, IO_5_77/DIFFIO_RX_R1N, IO_5_74/DIFFIO_RX_R2P, IO_5_75/DIFFIO_RX_R1P, IO_4_70/DIFFIO_TX_RX_B27P, IO_4_69/DIFFIO_TX_RX_B27N, IO_4_66/DIFFIO_TX_RX_B25N, IO_4_65/DIFFIO_TX_RX_B23P, IO_4_64/DIFFIO_TX_RX_B23N, IO_4_62/DIFFIO_TX_RX_B20P, IO_3_60/DIFFIO_TX_RX_B16P, IO_3_59/DIFFIO_TX_RX_B16N, IO_3_58/DIFFIO_TX_RX_B14P, IO_3_57/DIFFIO_TX_RX_B14N, IO_3_56/DIFFIO_TX_RX_B12P, IO_3_55/DIFFIO_TX_RX_B12N, IO_3_54/DIFFIO_TX_RX_B10N, IO_3_52/DIFFIO_TX_RX_B9P, IO_3_50/DIFFIO_TX_RX_B9N, IO_3_47/DIFFIO_TX_RX_B7P, IO_3_46/DIFFIO_TX_RX_B7N, IO_3_45/DIFFIO_TX_RX_B5P, IO_3_44/DIFFIO_TX_RX_B5N, IO_3_43/DIFFIO_TX_RX_B3P, IO_3_41/DIFFIO_TX_RX_B3N, IO_3_39/DIFFIO_TX_RX_B1P, IO_3_38/DIFFIO_TX_RX_B1N, IO_2_33/PLL_L_CLKOUTP/DIFFIO_RX_L27P, IO_2_32/PLL_L_CLKOUTN/DIFFIO_RX_L27N, IO_1B_25/DIFFIO_RX_L16P, IO_1B_24/DIFFIO_RX_L16N, IO_1B_22/DIFFIO_RX_L14P, IO_1B_21/DIFFIO_RX_L14N, IO_1A_14/ADC1IN8/DIFFIO_RX_L7P, IO_1A_13/ADC1IN7/DIFFIO_RX_L7N, IO_1A_12/ADC1IN6/DIFFIO_RX_L5P, IO_1A_11/ADC1IN5/DIFFIO_RX_L5N, IO_1A_10/ADC1IN4/DIFFIO_RX_L3P, IO_1A_8/ADC1IN3/DIFFIO_RX_L3N, IO_1A_7/ADC1IN2/DIFFIO_RX_L1P, IO_1A_6/ADC1IN1/DIFFIO_RX_L1N, VCC_ONE__1, VCC_ONE__108, VCC_ONE__109, VCC_ONE__115, VCC_ONE__144, VCC_ONE__36, VCC_ONE__37, VCC_ONE__51, VCC_ONE__72, VCC_ONE__73, VCCA6__2, VCCA5__71, VCCA4__143, VCCA3__107, VCCA2__34, VCCA1__35, VCCIO8__128, VCCIO8__139, VCCIO7__117, VCCIO6__103, VCCIO6__94, VCCIO5__82, VCCIO4__67, VCCIO3__40, VCCIO3__49, VCCIO2__31, VCCIO1B__23, VCCIO1A__9);

inout  Thermal;
inout  GND__142;

inout  GND__137;

inout  GND__133;

inout  GND__125;

inout  GND__116;

inout  GND__104;

inout  GND__95;

inout  GND__83;

inout  GND__68;

inout  GND__63;

inout  GND__53;

inout  GND__42;

inout  REFGND__4;

inout  ANAIN1__3;

inout  ADC_VREF__5;

inout  INPUT_ONLY_8_129/NCONFIG;
inout  IO_8_138/CONF_DONE/DIFFIO_RX_T24N;
inout  IO_8_136/NSTATUS/DIFFIO_RX_T24P;
inout  IO_8_134/CRC_ERROR/DIFFIO_RX_T22N;
inout  IO_8_126/BOOT_SEL;
inout  IO_8_122/DEV_OE/DIFFIO_RX_T18P;
inout  IO_8_121/DEV_CLRN/DIFFIO_RX_T16N;
inout  IO_1B_20/TDO/DIFFIO_RX_L12P;
inout  IO_1B_19/TDI/DIFFIO_RX_L12N;
inout  IO_1B_18/TCK/DIFFIO_RX_L11P;
inout  IO_1B_16/TMS/DIFFIO_RX_L11N;
inout  IO_1B_15/JTAGEN/DIFFIO_RX_L9P;
inout  IO_8_123/VREFB8N0;

inout  IO_7_112/VREFB7N0;

inout  IO_6_97/VREFB6N0;

inout  IO_5_80/VREFB5N0;

inout  IO_4_61/VREFB4N0;

inout  IO_3_48/VREFB3N0;

inout  IO_2_30/VREFB2N0;

inout  IO_1B_17/VREFB1N0;

inout  IO_6_98/DPCLK2/DIFFIO_RX_R26N;
inout  IO_6_96/DPCLK3/DIFFIO_RX_R26P;
inout  IO_6_91/CLK3N/DIFFIO_RX_R16N;
inout  IO_6_90/CLK3P/DIFFIO_RX_R16P;
inout  IO_6_89/CLK2N/DIFFIO_RX_R14N;
inout  IO_6_88/CLK2P/DIFFIO_RX_R14P;
inout  IO_2_29/CLK1P/DIFFIO_RX_L20P;
inout  IO_2_28/CLK1N/DIFFIO_RX_L20N;
inout  IO_2_27/CLK0P/DIFFIO_RX_L18P;
inout  IO_2_26/CLK0N/DIFFIO_RX_L18N;
inout  IO_8_120/DIFFIO_RX_T16P;
inout  IO_8_141/DIFFIO_RX_T26N;
inout  IO_8_140/DIFFIO_RX_T26P;
inout  IO_8_135/DIFFIO_RX_T23N;
inout  IO_8_132/DIFFIO_RX_T22P;
inout  IO_8_131/DIFFIO_RX_T20N;
inout  IO_8_130/DIFFIO_RX_T20P;
inout  IO_8_127/DIFFIO_RX_T19N;
inout  IO_8_124/DIFFIO_RX_T19P;
inout  IO_7_119/DIFFIO_RX_T10N;
inout  IO_7_118/DIFFIO_RX_T10P;
inout  IO_7_114/DIFFIO_RX_T6P;
inout  IO_7_113/DIFFIO_RX_T4N;
inout  IO_7_111/DIFFIO_RX_T1N;
inout  IO_7_110/DIFFIO_RX_T1P;
inout  IO_6_106/DIFFIO_RX_R33N;
inout  IO_6_105/DIFFIO_RX_R33P;
inout  IO_6_102/DIFFIO_RX_R28N;
inout  IO_6_101/DIFFIO_RX_R27N;
inout  IO_6_100/DIFFIO_RX_R28P;
inout  IO_6_99/DIFFIO_RX_R27P;
inout  IO_6_93/DIFFIO_RX_R18N;
inout  IO_6_92/DIFFIO_RX_R18P;
inout  IO_5_86/DIFFIO_RX_R11N;
inout  IO_5_87/DIFFIO_RX_R10N;
inout  IO_5_84/DIFFIO_RX_R11P;
inout  IO_5_85/DIFFIO_RX_R10P;
inout  IO_5_81/DIFFIO_RX_R7N;
inout  IO_5_78;

inout  IO_5_79/DIFFIO_RX_R7P;
inout  IO_5_76/DIFFIO_RX_R2N;
inout  IO_5_77/DIFFIO_RX_R1N;
inout  IO_5_74/DIFFIO_RX_R2P;
inout  IO_5_75/DIFFIO_RX_R1P;
inout  IO_4_70/DIFFIO_TX_RX_B27P;
inout  IO_4_69/DIFFIO_TX_RX_B27N;
inout  IO_4_66/DIFFIO_TX_RX_B25N;
inout  IO_4_65/DIFFIO_TX_RX_B23P;
inout  IO_4_64/DIFFIO_TX_RX_B23N;
inout  IO_4_62/DIFFIO_TX_RX_B20P;
inout  IO_3_60/DIFFIO_TX_RX_B16P;
inout  IO_3_59/DIFFIO_TX_RX_B16N;
inout  IO_3_58/DIFFIO_TX_RX_B14P;
inout  IO_3_57/DIFFIO_TX_RX_B14N;
inout  IO_3_56/DIFFIO_TX_RX_B12P;
inout  IO_3_55/DIFFIO_TX_RX_B12N;
inout  IO_3_54/DIFFIO_TX_RX_B10N;
inout  IO_3_52/DIFFIO_TX_RX_B9P;
inout  IO_3_50/DIFFIO_TX_RX_B9N;
inout  IO_3_47/DIFFIO_TX_RX_B7P;
inout  IO_3_46/DIFFIO_TX_RX_B7N;
inout  IO_3_45/DIFFIO_TX_RX_B5P;
inout  IO_3_44/DIFFIO_TX_RX_B5N;
inout  IO_3_43/DIFFIO_TX_RX_B3P;
inout  IO_3_41/DIFFIO_TX_RX_B3N;
inout  IO_3_39/DIFFIO_TX_RX_B1P;
inout  IO_3_38/DIFFIO_TX_RX_B1N;
inout  IO_2_33/PLL_L_CLKOUTP/DIFFIO_RX_L27P;
inout  IO_2_32/PLL_L_CLKOUTN/DIFFIO_RX_L27N;
inout  IO_1B_25/DIFFIO_RX_L16P;
inout  IO_1B_24/DIFFIO_RX_L16N;
inout  IO_1B_22/DIFFIO_RX_L14P;
inout  IO_1B_21/DIFFIO_RX_L14N;
inout  IO_1A_14/ADC1IN8/DIFFIO_RX_L7P;
inout  IO_1A_13/ADC1IN7/DIFFIO_RX_L7N;
inout  IO_1A_12/ADC1IN6/DIFFIO_RX_L5P;
inout  IO_1A_11/ADC1IN5/DIFFIO_RX_L5N;
inout  IO_1A_10/ADC1IN4/DIFFIO_RX_L3P;
inout  IO_1A_8/ADC1IN3/DIFFIO_RX_L3N;
inout  IO_1A_7/ADC1IN2/DIFFIO_RX_L1P;
inout  IO_1A_6/ADC1IN1/DIFFIO_RX_L1N;
inout  VCC_ONE__1;

inout  VCC_ONE__108;

inout  VCC_ONE__109;

inout  VCC_ONE__115;

inout  VCC_ONE__144;

inout  VCC_ONE__36;

inout  VCC_ONE__37;

inout  VCC_ONE__51;

inout  VCC_ONE__72;

inout  VCC_ONE__73;

inout  VCCA6__2;

inout  VCCA5__71;

inout  VCCA4__143;

inout  VCCA3__107;

inout  VCCA2__34;

inout  VCCA1__35;

inout  VCCIO8__128;

inout  VCCIO8__139;

inout  VCCIO7__117;

inout  VCCIO6__103;

inout  VCCIO6__94;

inout  VCCIO5__82;

inout  VCCIO4__67;

inout  VCCIO3__40;

inout  VCCIO3__49;

inout  VCCIO2__31;

inout  VCCIO1B__23;

inout  VCCIO1A__9;



endmodule
////////////////////////////////////////////////////////////////////////////////
